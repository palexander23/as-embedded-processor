//-----------------------------------------------------
// File Name        :   alucodes.sv
// Function         :   OPCODE Definitions
// Modified By      :   Peter Alexander
// Last rev. 24 Mar 2021
//-----------------------------------------------------

`define ACCI 2'b00
`define MACI 2'b01
`define BEQ  2'b10
`define BNE  2'b11
